library verilog;
use verilog.vl_types.all;
entity OPP_tb is
end OPP_tb;
